//-------------------------------------------------------------------------------------------------
// control center module 
// control initialization of all PEs 
//-------------------------------------------------------------------------------------------------

`timescale 1ns/1ps
import SystemVerilogCSP::*;
import dataformat::*;

module add
  #(parameter WIDTH = 5,
  parameter tot_num = 75,
  parameter tot_time = 3,
  parameter DATA_WIDTH = 20,
  parameter FL = 2,
  parameter BL = 2,
  parameter PACKDEALY = 1)

  ( input bit[WIDTH - 1:0] _index,
    input bit[WIDTH - 1:0] _mem_index,
    interface RouterToAdd_in,
    interface RouterToAdd_out,
    interface ccToAdd);

  int times[int];
  int sum[int];
  int pointer, i;
  bit flag = 0;
  bit[WIDTH - 1:0] index;
  bit[WIDTH - 1:0] mem_index;
  bit[DATA_WIDTH - 1:0] data_pass_memory;               
  bit[DATA_WIDTH - 1:0] data_pass_PE;                   

  always begin
      RouterToAdd_in.Receive(data_pass_PE);
      sum[data_pass_PE[DATA_WIDTH - 1:DATA_WIDTH-7]] += dataformater::unpackdata(data_pass_PE);
	  #PACKDEALY;
      times[data_pass_PE[DATA_WIDTH - 1:DATA_WIDTH-7]] += 1;
      #FL;
  end

  always begin
    wait(times[pointer] == tot_time);
    data_pass_memory = dataformater::packdata(index, mem_index, 0, sum[pointer]);
	#PACKDEALY;
    pointer = pointer + 1;
    RouterToAdd_out.Send(data_pass_memory);
    #BL;
  end

  always begin
    wait(pointer == tot_num);
    ccToAdd.Send(flag);
    #BL;
    ccToAdd.Receive(flag);
    #FL;
  end

  initial begin
    #0.1;
    pointer = 0;
    index = _index;
    mem_index = _mem_index;
    for(i = 0; i < tot_num; i = i + 1) begin
      times[i] = 0;
      sum[i] = 0;
    end
    ccToAdd.Receive(flag);
    #FL;
  end

endmodule
